library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package matrixmaker is
	type finalmatrix is array(0 to 7, 0 to 3) of unsigned (7 downto 0);
end package;