library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity main is
  port ();
end main;

architecture rtl of main is
begin
  -- codes
end rtl;
