
module PLL25 (
	clk_in_clk,
	clk_out_clk,
	clk_reset_reset);	

	input		clk_in_clk;
	output		clk_out_clk;
	input		clk_reset_reset;
endmodule
