-- library ieee;
-- use ieee.std_logic_1164.all;
-- use ieee.numeric_std.all;

-- package img_proc_pkg is
--         type img_arr is array(natural range <>) of std_logic_vector;
-- end package;

-- library ieee;
-- use ieee.std_logic_1164.all;
-- use ieee.numeric_std.all;
-- use work.img_proc_pkg.all;

-- entity img_proc is
--     port(
--         i_pixel : in img_arr(1)(3)
        
--     );
-- end img_proc;

-- architecture rtl of img_proc is

-- begin
    
-- end rtl;