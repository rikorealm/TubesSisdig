-- PLL25.vhd

-- Generated using ACDS version 23.1 993

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL25 is
	port (
		clk_in_clk      : in  std_logic := '0'; --    clk_in.clk
		clk_out_clk     : out std_logic;        --   clk_out.clk
		clk_reset_reset : in  std_logic := '0'  -- clk_reset.reset
	);
end entity PLL25;

architecture rtl of PLL25 is
	component PLL25_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component PLL25_altpll_0;

begin

	altpll_0 : component PLL25_altpll_0
		port map (
			clk                => clk_in_clk,      --       inclk_interface.clk
			reset              => clk_reset_reset, -- inclk_interface_reset.reset
			read               => open,            --             pll_slave.read
			write              => open,            --                      .write
			address            => open,            --                      .address
			readdata           => open,            --                      .readdata
			writedata          => open,            --                      .writedata
			c0                 => clk_out_clk,     --                    c0.clk
			scandone           => open,            --           (terminated)
			scandataout        => open,            --           (terminated)
			areset             => '0',             --           (terminated)
			locked             => open,            --           (terminated)
			phasedone          => open,            --           (terminated)
			phasecounterselect => "0000",          --           (terminated)
			phaseupdown        => '0',             --           (terminated)
			phasestep          => '0',             --           (terminated)
			scanclk            => '0',             --           (terminated)
			scanclkena         => '0',             --           (terminated)
			scandata           => '0',             --           (terminated)
			configupdate       => '0'              --           (terminated)
		);

end architecture rtl; -- of PLL25
